`timescale 1ns/1ps
// 2000 ciclos para responder

module tb_fpu;
    reg clk;
    reg reset;

    initial begin
        $dumpfile("tb_fpu.vcd");
        $dumpvars(0,tb_fpu);
    end

    always #1 clk = !clk;

    reg [31:0] A, B;
    reg [1:0] op;
    reg start;
    wire [31:0] R;
    wire done;

    fpu fpu (clk, reset, A, B, R, op, start, done);

    initial begin
        #1;
        reset = 0;
        start = 1;

        op = 2'b00;

        A = 32'b00111111101000000000000000000000;
        B = 32'b00111111110000000000000000000000;
        // 1,25 + 1,5

        #200;

        start = 0;
        #2;
        start = 1;

        A = 32'b01000010001010101010111000010100;
        B = 32'b01000010000100001100110011001101;
        // possible roundind error
        // 42,67 + 36,2 = 78,87
        #200;

        start = 0;
        #2;
        start = 1;

        A = 32'b00111011101000111101011100001010;
        B = 32'b00111110000011110101110000101001;
        // 0,005 + 0,14 = 0,145
        #200;

        start = 0;
        #2;
        start = 1;

        A = 32'b00111110100010100011110101110001;
        B = 32'b01000000100111110101110000101001;
        // 0,27 + 4,98 = 5,25

        #200;

        start = 0;
        #2;
        start = 1;

        A = 32'b01000000111000000000000000000000;
        B = 32'b01000000111110000000000000000000;
        // 7,0 + 7,75 = 14,75

        #200;
        start = 0;
        #2;
        start = 1;

        A = 32'b01000001110011000000000000000000;
        B = 32'b01000001111011000000000000000000;
        // 25,5 + 29,5 = 55

        #200;
        start = 0;
        #2;
        start = 1;

        A = 32'b00111111110000000000000000000000;
        B = 32'b00000000000000000000000000000000;
        // 1,5 + 0 = 1,5

        #200;
        start = 0;
        #2;
        start = 1;

        A = 32'b11000000001100000000000000000000;
        B = 32'b11000000010100000000000000000000;
        // -2,75 - 3,25 = -6

        #200;
        start = 0;
        #2;
        start = 1;

        A = 32'b10111111010000000000000000000000;
        B = 32'b00111110100000000000000000000000;
        // -0,75 + 0,25 = -0,5
        #200;

        start = 0;
        op = 2'b10;
        #2;
        start = 1;

        A = 32'b01000000001000000000000000000000;
        B = 32'b01000000100110000000000000000000;
        // 2.5 * 4,75 = 11,875
        #200;

        start = 0;
        #2;
        start = 1;

        A = 32'b10111110000000000000000000000000;
        B = 32'b10111110111000000000000000000000;
        // -1,125 * -0.4375 = 0.4921875
        #200;

        start = 0;
        #2;
        start = 1;

        A = 32'b00111111010101000000000000000000;
        B = 32'b11000001010101000000000000000000;
        // 0.828125 * -13.25 = -10,97265625
        #200;

        $finish;
    end

    initial begin
        $monitor("A = %b | B = %b | R = %b", A, B, R);
    end

endmodule