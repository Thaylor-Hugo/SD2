// memoria rom para multiplicacao de numeros de 5 bits e saida de 10

module rom (
    input [9:0] endereco,
    output [9:0] resultado
);

reg [9:0] rom [1023:0];
integer i, j;

initial begin
    rom[0] = 0;
    rom[1] = 0;
    rom[2] = 0;
    rom[3] = 0;
    rom[4] = 0;
    rom[5] = 0;
    rom[6] = 0;
    rom[7] = 0;
    rom[8] = 0;
    rom[9] = 0;
    rom[10] = 0;
    rom[11] = 0;
    rom[12] = 0;
    rom[13] = 0;
    rom[14] = 0;
    rom[15] = 0;
    rom[16] = 0;
    rom[17] = 0;
    rom[18] = 0;
    rom[19] = 0;
    rom[20] = 0;
    rom[21] = 0;
    rom[22] = 0;
    rom[23] = 0;
    rom[24] = 0;
    rom[25] = 0;
    rom[26] = 0;
    rom[27] = 0;
    rom[28] = 0;
    rom[29] = 0;
    rom[30] = 0;
    rom[31] = 0;
    rom[32] = 0;
    rom[33] = 1;
    rom[34] = 2;
    rom[35] = 3;
    rom[36] = 4;
    rom[37] = 5;
    rom[38] = 6;
    rom[39] = 7;
    rom[40] = 8;
    rom[41] = 9;
    rom[42] = 10;
    rom[43] = 11;
    rom[44] = 12;
    rom[45] = 13;
    rom[46] = 14;
    rom[47] = 15;
    rom[48] = 16;
    rom[49] = 17;
    rom[50] = 18;
    rom[51] = 19;
    rom[52] = 20;
    rom[53] = 21;
    rom[54] = 22;
    rom[55] = 23;
    rom[56] = 24;
    rom[57] = 25;
    rom[58] = 26;
    rom[59] = 27;
    rom[60] = 28;
    rom[61] = 29;
    rom[62] = 30;
    rom[63] = 31;
    rom[64] = 0;
    rom[65] = 2;
    rom[66] = 4;
    rom[67] = 6;
    rom[68] = 8;
    rom[69] = 10;
    rom[70] = 12;
    rom[71] = 14;
    rom[72] = 16;
    rom[73] = 18;
    rom[74] = 20;
    rom[75] = 22;
    rom[76] = 24;
    rom[77] = 26;
    rom[78] = 28;
    rom[79] = 30;
    rom[80] = 32;
    rom[81] = 34;
    rom[82] = 36;
    rom[83] = 38;
    rom[84] = 40;
    rom[85] = 42;
    rom[86] = 44;
    rom[87] = 46;
    rom[88] = 48;
    rom[89] = 50;
    rom[90] = 52;
    rom[91] = 54;
    rom[92] = 56;
    rom[93] = 58;
    rom[94] = 60;
    rom[95] = 62;
    rom[96] = 0;
    rom[97] = 3;
    rom[98] = 6;
    rom[99] = 9;
    rom[100] = 12;
    rom[101] = 15;
    rom[102] = 18;
    rom[103] = 21;
    rom[104] = 24;
    rom[105] = 27;
    rom[106] = 30;
    rom[107] = 33;
    rom[108] = 36;
    rom[109] = 39;
    rom[110] = 42;
    rom[111] = 45;
    rom[112] = 48;
    rom[113] = 51;
    rom[114] = 54;
    rom[115] = 57;
    rom[116] = 60;
    rom[117] = 63;
    rom[118] = 66;
    rom[119] = 69;
    rom[120] = 72;
    rom[121] = 75;
    rom[122] = 78;
    rom[123] = 81;
    rom[124] = 84;
    rom[125] = 87;
    rom[126] = 90;
    rom[127] = 93;
    rom[128] = 0;
    rom[129] = 4;
    rom[130] = 8;
    rom[131] = 12;
    rom[132] = 16;
    rom[133] = 20;
    rom[134] = 24;
    rom[135] = 28;
    rom[136] = 32;
    rom[137] = 36;
    rom[138] = 40;
    rom[139] = 44;
    rom[140] = 48;
    rom[141] = 52;
    rom[142] = 56;
    rom[143] = 60;
    rom[144] = 64;
    rom[145] = 68;
    rom[146] = 72;
    rom[147] = 76;
    rom[148] = 80;
    rom[149] = 84;
    rom[150] = 88;
    rom[151] = 92;
    rom[152] = 96;
    rom[153] = 100;
    rom[154] = 104;
    rom[155] = 108;
    rom[156] = 112;
    rom[157] = 116;
    rom[158] = 120;
    rom[159] = 124;
    rom[160] = 0;
    rom[161] = 5;
    rom[162] = 10;
    rom[163] = 15;
    rom[164] = 20;
    rom[165] = 25;
    rom[166] = 30;
    rom[167] = 35;
    rom[168] = 40;
    rom[169] = 45;
    rom[170] = 50;
    rom[171] = 55;
    rom[172] = 60;
    rom[173] = 65;
    rom[174] = 70;
    rom[175] = 75;
    rom[176] = 80;
    rom[177] = 85;
    rom[178] = 90;
    rom[179] = 95;
    rom[180] = 100;
    rom[181] = 105;
    rom[182] = 110;
    rom[183] = 115;
    rom[184] = 120;
    rom[185] = 125;
    rom[186] = 130;
    rom[187] = 135;
    rom[188] = 140;
    rom[189] = 145;
    rom[190] = 150;
    rom[191] = 155;
    rom[192] = 0;
    rom[193] = 6;
    rom[194] = 12;
    rom[195] = 18;
    rom[196] = 24;
    rom[197] = 30;
    rom[198] = 36;
    rom[199] = 42;
    rom[200] = 48;
    rom[201] = 54;
    rom[202] = 60;
    rom[203] = 66;
    rom[204] = 72;
    rom[205] = 78;
    rom[206] = 84;
    rom[207] = 90;
    rom[208] = 96;
    rom[209] = 102;
    rom[210] = 108;
    rom[211] = 114;
    rom[212] = 120;
    rom[213] = 126;
    rom[214] = 132;
    rom[215] = 138;
    rom[216] = 144;
    rom[217] = 150;
    rom[218] = 156;
    rom[219] = 162;
    rom[220] = 168;
    rom[221] = 174;
    rom[222] = 180;
    rom[223] = 186;
    rom[224] = 0;
    rom[225] = 7;
    rom[226] = 14;
    rom[227] = 21;
    rom[228] = 28;
    rom[229] = 35;
    rom[230] = 42;
    rom[231] = 49;
    rom[232] = 56;
    rom[233] = 63;
    rom[234] = 70;
    rom[235] = 77;
    rom[236] = 84;
    rom[237] = 91;
    rom[238] = 98;
    rom[239] = 105;
    rom[240] = 112;
    rom[241] = 119;
    rom[242] = 126;
    rom[243] = 133;
    rom[244] = 140;
    rom[245] = 147;
    rom[246] = 154;
    rom[247] = 161;
    rom[248] = 168;
    rom[249] = 175;
    rom[250] = 182;
    rom[251] = 189;
    rom[252] = 196;
    rom[253] = 203;
    rom[254] = 210;
    rom[255] = 217;
    rom[256] = 0;
    rom[257] = 8;
    rom[258] = 16;
    rom[259] = 24;
    rom[260] = 32;
    rom[261] = 40;
    rom[262] = 48;
    rom[263] = 56;
    rom[264] = 64;
    rom[265] = 72;
    rom[266] = 80;
    rom[267] = 88;
    rom[268] = 96;
    rom[269] = 104;
    rom[270] = 112;
    rom[271] = 120;
    rom[272] = 128;
    rom[273] = 136;
    rom[274] = 144;
    rom[275] = 152;
    rom[276] = 160;
    rom[277] = 168;
    rom[278] = 176;
    rom[279] = 184;
    rom[280] = 192;
    rom[281] = 200;
    rom[282] = 208;
    rom[283] = 216;
    rom[284] = 224;
    rom[285] = 232;
    rom[286] = 240;
    rom[287] = 248;
    rom[288] = 0;
    rom[289] = 9;
    rom[290] = 18;
    rom[291] = 27;
    rom[292] = 36;
    rom[293] = 45;
    rom[294] = 54;
    rom[295] = 63;
    rom[296] = 72;
    rom[297] = 81;
    rom[298] = 90;
    rom[299] = 99;
    rom[300] = 108;
    rom[301] = 117;
    rom[302] = 126;
    rom[303] = 135;
    rom[304] = 144;
    rom[305] = 153;
    rom[306] = 162;
    rom[307] = 171;
    rom[308] = 180;
    rom[309] = 189;
    rom[310] = 198;
    rom[311] = 207;
    rom[312] = 216;
    rom[313] = 225;
    rom[314] = 234;
    rom[315] = 243;
    rom[316] = 252;
    rom[317] = 261;
    rom[318] = 270;
    rom[319] = 279;
    rom[320] = 0;
    rom[321] = 10;
    rom[322] = 20;
    rom[323] = 30;
    rom[324] = 40;
    rom[325] = 50;
    rom[326] = 60;
    rom[327] = 70;
    rom[328] = 80;
    rom[329] = 90;
    rom[330] = 100;
    rom[331] = 110;
    rom[332] = 120;
    rom[333] = 130;
    rom[334] = 140;
    rom[335] = 150;
    rom[336] = 160;
    rom[337] = 170;
    rom[338] = 180;
    rom[339] = 190;
    rom[340] = 200;
    rom[341] = 210;
    rom[342] = 220;
    rom[343] = 230;
    rom[344] = 240;
    rom[345] = 250;
    rom[346] = 260;
    rom[347] = 270;
    rom[348] = 280;
    rom[349] = 290;
    rom[350] = 300;
    rom[351] = 310;
    rom[352] = 0;
    rom[353] = 11;
    rom[354] = 22;
    rom[355] = 33;
    rom[356] = 44;
    rom[357] = 55;
    rom[358] = 66;
    rom[359] = 77;
    rom[360] = 88;
    rom[361] = 99;
    rom[362] = 110;
    rom[363] = 121;
    rom[364] = 132;
    rom[365] = 143;
    rom[366] = 154;
    rom[367] = 165;
    rom[368] = 176;
    rom[369] = 187;
    rom[370] = 198;
    rom[371] = 209;
    rom[372] = 220;
    rom[373] = 231;
    rom[374] = 242;
    rom[375] = 253;
    rom[376] = 264;
    rom[377] = 275;
    rom[378] = 286;
    rom[379] = 297;
    rom[380] = 308;
    rom[381] = 319;
    rom[382] = 330;
    rom[383] = 341;
    rom[384] = 0;
    rom[385] = 12;
    rom[386] = 24;
    rom[387] = 36;
    rom[388] = 48;
    rom[389] = 60;
    rom[390] = 72;
    rom[391] = 84;
    rom[392] = 96;
    rom[393] = 108;
    rom[394] = 120;
    rom[395] = 132;
    rom[396] = 144;
    rom[397] = 156;
    rom[398] = 168;
    rom[399] = 180;
    rom[400] = 192;
    rom[401] = 204;
    rom[402] = 216;
    rom[403] = 228;
    rom[404] = 240;
    rom[405] = 252;
    rom[406] = 264;
    rom[407] = 276;
    rom[408] = 288;
    rom[409] = 300;
    rom[410] = 312;
    rom[411] = 324;
    rom[412] = 336;
    rom[413] = 348;
    rom[414] = 360;
    rom[415] = 372;
    rom[416] = 0;
    rom[417] = 13;
    rom[418] = 26;
    rom[419] = 39;
    rom[420] = 52;
    rom[421] = 65;
    rom[422] = 78;
    rom[423] = 91;
    rom[424] = 104;
    rom[425] = 117;
    rom[426] = 130;
    rom[427] = 143;
    rom[428] = 156;
    rom[429] = 169;
    rom[430] = 182;
    rom[431] = 195;
    rom[432] = 208;
    rom[433] = 221;
    rom[434] = 234;
    rom[435] = 247;
    rom[436] = 260;
    rom[437] = 273;
    rom[438] = 286;
    rom[439] = 299;
    rom[440] = 312;
    rom[441] = 325;
    rom[442] = 338;
    rom[443] = 351;
    rom[444] = 364;
    rom[445] = 377;
    rom[446] = 390;
    rom[447] = 403;
    rom[448] = 0;
    rom[449] = 14;
    rom[450] = 28;
    rom[451] = 42;
    rom[452] = 56;
    rom[453] = 70;
    rom[454] = 84;
    rom[455] = 98;
    rom[456] = 112;
    rom[457] = 126;
    rom[458] = 140;
    rom[459] = 154;
    rom[460] = 168;
    rom[461] = 182;
    rom[462] = 196;
    rom[463] = 210;
    rom[464] = 224;
    rom[465] = 238;
    rom[466] = 252;
    rom[467] = 266;
    rom[468] = 280;
    rom[469] = 294;
    rom[470] = 308;
    rom[471] = 322;
    rom[472] = 336;
    rom[473] = 350;
    rom[474] = 364;
    rom[475] = 378;
    rom[476] = 392;
    rom[477] = 406;
    rom[478] = 420;
    rom[479] = 434;
    rom[480] = 0;
    rom[481] = 15;
    rom[482] = 30;
    rom[483] = 45;
    rom[484] = 60;
    rom[485] = 75;
    rom[486] = 90;
    rom[487] = 105;
    rom[488] = 120;
    rom[489] = 135;
    rom[490] = 150;
    rom[491] = 165;
    rom[492] = 180;
    rom[493] = 195;
    rom[494] = 210;
    rom[495] = 225;
    rom[496] = 240;
    rom[497] = 255;
    rom[498] = 270;
    rom[499] = 285;
    rom[500] = 300;
    rom[501] = 315;
    rom[502] = 330;
    rom[503] = 345;
    rom[504] = 360;
    rom[505] = 375;
    rom[506] = 390;
    rom[507] = 405;
    rom[508] = 420;
    rom[509] = 435;
    rom[510] = 450;
    rom[511] = 465;
    rom[512] = 0;
    rom[513] = 16;
    rom[514] = 32;
    rom[515] = 48;
    rom[516] = 64;
    rom[517] = 80;
    rom[518] = 96;
    rom[519] = 112;
    rom[520] = 128;
    rom[521] = 144;
    rom[522] = 160;
    rom[523] = 176;
    rom[524] = 192;
    rom[525] = 208;
    rom[526] = 224;
    rom[527] = 240;
    rom[528] = 256;
    rom[529] = 272;
    rom[530] = 288;
    rom[531] = 304;
    rom[532] = 320;
    rom[533] = 336;
    rom[534] = 352;
    rom[535] = 368;
    rom[536] = 384;
    rom[537] = 400;
    rom[538] = 416;
    rom[539] = 432;
    rom[540] = 448;
    rom[541] = 464;
    rom[542] = 480;
    rom[543] = 496;
    rom[544] = 0;
    rom[545] = 17;
    rom[546] = 34;
    rom[547] = 51;
    rom[548] = 68;
    rom[549] = 85;
    rom[550] = 102;
    rom[551] = 119;
    rom[552] = 136;
    rom[553] = 153;
    rom[554] = 170;
    rom[555] = 187;
    rom[556] = 204;
    rom[557] = 221;
    rom[558] = 238;
    rom[559] = 255;
    rom[560] = 272;
    rom[561] = 289;
    rom[562] = 306;
    rom[563] = 323;
    rom[564] = 340;
    rom[565] = 357;
    rom[566] = 374;
    rom[567] = 391;
    rom[568] = 408;
    rom[569] = 425;
    rom[570] = 442;
    rom[571] = 459;
    rom[572] = 476;
    rom[573] = 493;
    rom[574] = 510;
    rom[575] = 527;
    rom[576] = 0;
    rom[577] = 18;
    rom[578] = 36;
    rom[579] = 54;
    rom[580] = 72;
    rom[581] = 90;
    rom[582] = 108;
    rom[583] = 126;
    rom[584] = 144;
    rom[585] = 162;
    rom[586] = 180;
    rom[587] = 198;
    rom[588] = 216;
    rom[589] = 234;
    rom[590] = 252;
    rom[591] = 270;
    rom[592] = 288;
    rom[593] = 306;
    rom[594] = 324;
    rom[595] = 342;
    rom[596] = 360;
    rom[597] = 378;
    rom[598] = 396;
    rom[599] = 414;
    rom[600] = 432;
    rom[601] = 450;
    rom[602] = 468;
    rom[603] = 486;
    rom[604] = 504;
    rom[605] = 522;
    rom[606] = 540;
    rom[607] = 558;
    rom[608] = 0;
    rom[609] = 19;
    rom[610] = 38;
    rom[611] = 57;
    rom[612] = 76;
    rom[613] = 95;
    rom[614] = 114;
    rom[615] = 133;
    rom[616] = 152;
    rom[617] = 171;
    rom[618] = 190;
    rom[619] = 209;
    rom[620] = 228;
    rom[621] = 247;
    rom[622] = 266;
    rom[623] = 285;
    rom[624] = 304;
    rom[625] = 323;
    rom[626] = 342;
    rom[627] = 361;
    rom[628] = 380;
    rom[629] = 399;
    rom[630] = 418;
    rom[631] = 437;
    rom[632] = 456;
    rom[633] = 475;
    rom[634] = 494;
    rom[635] = 513;
    rom[636] = 532;
    rom[637] = 551;
    rom[638] = 570;
    rom[639] = 589;
    rom[640] = 0;
    rom[641] = 20;
    rom[642] = 40;
    rom[643] = 60;
    rom[644] = 80;
    rom[645] = 100;
    rom[646] = 120;
    rom[647] = 140;
    rom[648] = 160;
    rom[649] = 180;
    rom[650] = 200;
    rom[651] = 220;
    rom[652] = 240;
    rom[653] = 260;
    rom[654] = 280;
    rom[655] = 300;
    rom[656] = 320;
    rom[657] = 340;
    rom[658] = 360;
    rom[659] = 380;
    rom[660] = 400;
    rom[661] = 420;
    rom[662] = 440;
    rom[663] = 460;
    rom[664] = 480;
    rom[665] = 500;
    rom[666] = 520;
    rom[667] = 540;
    rom[668] = 560;
    rom[669] = 580;
    rom[670] = 600;
    rom[671] = 620;
    rom[672] = 0;
    rom[673] = 21;
    rom[674] = 42;
    rom[675] = 63;
    rom[676] = 84;
    rom[677] = 105;
    rom[678] = 126;
    rom[679] = 147;
    rom[680] = 168;
    rom[681] = 189;
    rom[682] = 210;
    rom[683] = 231;
    rom[684] = 252;
    rom[685] = 273;
    rom[686] = 294;
    rom[687] = 315;
    rom[688] = 336;
    rom[689] = 357;
    rom[690] = 378;
    rom[691] = 399;
    rom[692] = 420;
    rom[693] = 441;
    rom[694] = 462;
    rom[695] = 483;
    rom[696] = 504;
    rom[697] = 525;
    rom[698] = 546;
    rom[699] = 567;
    rom[700] = 588;
    rom[701] = 609;
    rom[702] = 630;
    rom[703] = 651;
    rom[704] = 0;
    rom[705] = 22;
    rom[706] = 44;
    rom[707] = 66;
    rom[708] = 88;
    rom[709] = 110;
    rom[710] = 132;
    rom[711] = 154;
    rom[712] = 176;
    rom[713] = 198;
    rom[714] = 220;
    rom[715] = 242;
    rom[716] = 264;
    rom[717] = 286;
    rom[718] = 308;
    rom[719] = 330;
    rom[720] = 352;
    rom[721] = 374;
    rom[722] = 396;
    rom[723] = 418;
    rom[724] = 440;
    rom[725] = 462;
    rom[726] = 484;
    rom[727] = 506;
    rom[728] = 528;
    rom[729] = 550;
    rom[730] = 572;
    rom[731] = 594;
    rom[732] = 616;
    rom[733] = 638;
    rom[734] = 660;
    rom[735] = 682;
    rom[736] = 0;
    rom[737] = 23;
    rom[738] = 46;
    rom[739] = 69;
    rom[740] = 92;
    rom[741] = 115;
    rom[742] = 138;
    rom[743] = 161;
    rom[744] = 184;
    rom[745] = 207;
    rom[746] = 230;
    rom[747] = 253;
    rom[748] = 276;
    rom[749] = 299;
    rom[750] = 322;
    rom[751] = 345;
    rom[752] = 368;
    rom[753] = 391;
    rom[754] = 414;
    rom[755] = 437;
    rom[756] = 460;
    rom[757] = 483;
    rom[758] = 506;
    rom[759] = 529;
    rom[760] = 552;
    rom[761] = 575;
    rom[762] = 598;
    rom[763] = 621;
    rom[764] = 644;
    rom[765] = 667;
    rom[766] = 690;
    rom[767] = 713;
    rom[768] = 0;
    rom[769] = 24;
    rom[770] = 48;
    rom[771] = 72;
    rom[772] = 96;
    rom[773] = 120;
    rom[774] = 144;
    rom[775] = 168;
    rom[776] = 192;
    rom[777] = 216;
    rom[778] = 240;
    rom[779] = 264;
    rom[780] = 288;
    rom[781] = 312;
    rom[782] = 336;
    rom[783] = 360;
    rom[784] = 384;
    rom[785] = 408;
    rom[786] = 432;
    rom[787] = 456;
    rom[788] = 480;
    rom[789] = 504;
    rom[790] = 528;
    rom[791] = 552;
    rom[792] = 576;
    rom[793] = 600;
    rom[794] = 624;
    rom[795] = 648;
    rom[796] = 672;
    rom[797] = 696;
    rom[798] = 720;
    rom[799] = 744;
    rom[800] = 0;
    rom[801] = 25;
    rom[802] = 50;
    rom[803] = 75;
    rom[804] = 100;
    rom[805] = 125;
    rom[806] = 150;
    rom[807] = 175;
    rom[808] = 200;
    rom[809] = 225;
    rom[810] = 250;
    rom[811] = 275;
    rom[812] = 300;
    rom[813] = 325;
    rom[814] = 350;
    rom[815] = 375;
    rom[816] = 400;
    rom[817] = 425;
    rom[818] = 450;
    rom[819] = 475;
    rom[820] = 500;
    rom[821] = 525;
    rom[822] = 550;
    rom[823] = 575;
    rom[824] = 600;
    rom[825] = 625;
    rom[826] = 650;
    rom[827] = 675;
    rom[828] = 700;
    rom[829] = 725;
    rom[830] = 750;
    rom[831] = 775;
    rom[832] = 0;
    rom[833] = 26;
    rom[834] = 52;
    rom[835] = 78;
    rom[836] = 104;
    rom[837] = 130;
    rom[838] = 156;
    rom[839] = 182;
    rom[840] = 208;
    rom[841] = 234;
    rom[842] = 260;
    rom[843] = 286;
    rom[844] = 312;
    rom[845] = 338;
    rom[846] = 364;
    rom[847] = 390;
    rom[848] = 416;
    rom[849] = 442;
    rom[850] = 468;
    rom[851] = 494;
    rom[852] = 520;
    rom[853] = 546;
    rom[854] = 572;
    rom[855] = 598;
    rom[856] = 624;
    rom[857] = 650;
    rom[858] = 676;
    rom[859] = 702;
    rom[860] = 728;
    rom[861] = 754;
    rom[862] = 780;
    rom[863] = 806;
    rom[864] = 0;
    rom[865] = 27;
    rom[866] = 54;
    rom[867] = 81;
    rom[868] = 108;
    rom[869] = 135;
    rom[870] = 162;
    rom[871] = 189;
    rom[872] = 216;
    rom[873] = 243;
    rom[874] = 270;
    rom[875] = 297;
    rom[876] = 324;
    rom[877] = 351;
    rom[878] = 378;
    rom[879] = 405;
    rom[880] = 432;
    rom[881] = 459;
    rom[882] = 486;
    rom[883] = 513;
    rom[884] = 540;
    rom[885] = 567;
    rom[886] = 594;
    rom[887] = 621;
    rom[888] = 648;
    rom[889] = 675;
    rom[890] = 702;
    rom[891] = 729;
    rom[892] = 756;
    rom[893] = 783;
    rom[894] = 810;
    rom[895] = 837;
    rom[896] = 0;
    rom[897] = 28;
    rom[898] = 56;
    rom[899] = 84;
    rom[900] = 112;
    rom[901] = 140;
    rom[902] = 168;
    rom[903] = 196;
    rom[904] = 224;
    rom[905] = 252;
    rom[906] = 280;
    rom[907] = 308;
    rom[908] = 336;
    rom[909] = 364;
    rom[910] = 392;
    rom[911] = 420;
    rom[912] = 448;
    rom[913] = 476;
    rom[914] = 504;
    rom[915] = 532;
    rom[916] = 560;
    rom[917] = 588;
    rom[918] = 616;
    rom[919] = 644;
    rom[920] = 672;
    rom[921] = 700;
    rom[922] = 728;
    rom[923] = 756;
    rom[924] = 784;
    rom[925] = 812;
    rom[926] = 840;
    rom[927] = 868;
    rom[928] = 0;
    rom[929] = 29;
    rom[930] = 58;
    rom[931] = 87;
    rom[932] = 116;
    rom[933] = 145;
    rom[934] = 174;
    rom[935] = 203;
    rom[936] = 232;
    rom[937] = 261;
    rom[938] = 290;
    rom[939] = 319;
    rom[940] = 348;
    rom[941] = 377;
    rom[942] = 406;
    rom[943] = 435;
    rom[944] = 464;
    rom[945] = 493;
    rom[946] = 522;
    rom[947] = 551;
    rom[948] = 580;
    rom[949] = 609;
    rom[950] = 638;
    rom[951] = 667;
    rom[952] = 696;
    rom[953] = 725;
    rom[954] = 754;
    rom[955] = 783;
    rom[956] = 812;
    rom[957] = 841;
    rom[958] = 870;
    rom[959] = 899;
    rom[960] = 0;
    rom[961] = 30;
    rom[962] = 60;
    rom[963] = 90;
    rom[964] = 120;
    rom[965] = 150;
    rom[966] = 180;
    rom[967] = 210;
    rom[968] = 240;
    rom[969] = 270;
    rom[970] = 300;
    rom[971] = 330;
    rom[972] = 360;
    rom[973] = 390;
    rom[974] = 420;
    rom[975] = 450;
    rom[976] = 480;
    rom[977] = 510;
    rom[978] = 540;
    rom[979] = 570;
    rom[980] = 600;
    rom[981] = 630;
    rom[982] = 660;
    rom[983] = 690;
    rom[984] = 720;
    rom[985] = 750;
    rom[986] = 780;
    rom[987] = 810;
    rom[988] = 840;
    rom[989] = 870;
    rom[990] = 900;
    rom[991] = 930;
    rom[992] = 0;
    rom[993] = 31;
    rom[994] = 62;
    rom[995] = 93;
    rom[996] = 124;
    rom[997] = 155;
    rom[998] = 186;
    rom[999] = 217;
    rom[1000] = 248;
    rom[1001] = 279;
    rom[1002] = 310;
    rom[1003] = 341;
    rom[1004] = 372;
    rom[1005] = 403;
    rom[1006] = 434;
    rom[1007] = 465;
    rom[1008] = 496;
    rom[1009] = 527;
    rom[1010] = 558;
    rom[1011] = 589;
    rom[1012] = 620;
    rom[1013] = 651;
    rom[1014] = 682;
    rom[1015] = 713;
    rom[1016] = 744;
    rom[1017] = 775;
    rom[1018] = 806;
    rom[1019] = 837;
    rom[1020] = 868;
    rom[1021] = 899;
    rom[1022] = 930;
    rom[1023] = 961;
end

assign resultado = rom[endereco];
    
endmodule