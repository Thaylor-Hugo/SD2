// Grupo 5
// Nomes:
// Thaylor Hugo - 13684425 
// Felipe Soria - 13864287
// Alejandro Larrea - 13791522  

// ULA em complemento de 2
module somador (
    input [7:0] a,
    input [7:0] b,
    output [7:0] result
);

assign result = a + b;

endmodule
